//===============================================================
// File Name        : mvt_clk_interface
// Description      :
// Name             : zhangjunxiao
// File Created     : 01/06/2025 @ 05:18 PM
// Copyright        :
//===============================================================
// NOTE: Please Don't Remove Any Comments or //--- Given Below
//===============================================================

//---------------------------------------------------------------
// Interface: mvt_clk_interface
// 
//---------------------------------------------------------------

interface mvt_clk_interface ;
 //------------------------------------------
 // Signal Instantiation
 //------------------------------------------
endinterface: mvt_clk_interface

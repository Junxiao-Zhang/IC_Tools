module gddr6_checker (
    input        CLK,
    input        CLKB,
    input        WCLK0,
    input        WCLK0B,
    input        WCLK1,
    input        WCLK1B,
    input        CKEB,
    input        CABIB,
    input [10:0] CA,
    input [15:0] DQ,
    input [ 1:0] DBIB,
    input [ 1:0] EDC,
    input        RESETB

);

endmodule
